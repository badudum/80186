

module execUnit();


endmodule

