

module biu ()

endmodule