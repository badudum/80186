

`timescale 1ns/1ns
module ALU()
//TODO : CREATE THIS MODULE

endmodule 